`timescale 1ns / 1ps
module alto_io_controller (
	input clk_i,
	input rst_i,
	
	output sck_o,
	output mosi_o,
	input miso_i,
	output ss_o
);


endmodule
